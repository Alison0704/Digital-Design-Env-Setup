module top_module(
  // ports
);
  // TODO: implement
endmodule
