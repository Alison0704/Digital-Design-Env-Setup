module top_module(
  // TODO: implement ports
);
  // TODO: implement
endmodule
