library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity top_module is
    Port (
           -- // TODO:  define the ports
    );
end top_module;

architecture Behavioral of top_module is
    -- Declare internal signals here
begin
    -- // TODO: implement the processes
end Behavioral;